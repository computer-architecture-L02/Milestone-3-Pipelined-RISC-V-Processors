module alu()
endmodule
